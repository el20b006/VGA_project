-------------------------------------------------------------------------------
--                                                                      
--                        VGA Controller VHDL Project
--  
-------------------------------------------------------------------------------
--                                                                      
-- ENTITY:         VGA_ctrl_top
--
-- FILENAME:       VGA_ctrl_top_struc_cfg.vhd
-- 
-- ARCHITECTURE:   struc
-- 
-- ENGINEER:       Sarah Fr�ler
--
-- DATE:           16. January 2023
--
-- VERSION:        1.0
--
-------------------------------------------------------------------------------
--                                                                      
-- DESCRIPTION:    This is the configuration for the entity VGA_ctrl_top and 
--                 the architecture struc.
--
--
-------------------------------------------------------------------------------
--
-- REFERENCES:     (none)
--
-------------------------------------------------------------------------------
--                                                                      
-- PACKAGES:       std_logic_1164 (IEEE library)
--
-------------------------------------------------------------------------------
--                                                                      
-- CHANGES:        Version 1.0
--
-------------------------------------------------------------------------------

configuration VGA_ctrl_top_struc_cfg of VGA_ctrl_top is
  for struc      -- architecture struc is used for entity VGA top
  end for;
end VGA_ctrl_top_struc_cfg;
